module BC82AMDD_CPLD1
 (
 input  Test1,
 input  test2,
 
 )
  
  
  
endmodule
